.MODEL 1N4148W D  ( IS=10.4n RS=51.5m BV=75.0 IBV=1.00u
+ CJO=2.00p  M=0.333 N=2.07 TT=5.76n )
V1 0 in DC 5
R1 in 1 11.72
R2 1 2 220
D1 2 0 1N4148W